r1 1 0 1
i1 0 1 10
r2 1 2 100
r3 2 3 100
r4 3 4 100
r5 4 0 100
