i1 0 1 2
r1 1 2 1
r2 2 0 1
x1 3 4 1 2 10
r3 3 0 1
r4 4 0 1
